`timescale 1ns / 1ps
module LUT_bias ( Iin, Out);


input  [7:0] Iin;
output reg [31:0] Out;

always @ *//( posedge En )
begin 
case (Iin)

8'b10000000 : Out =32'b00000000000000000000000000000000;
8'b10000001 : Out =32'b00000000000000000000000000000000;
8'b10000010 : Out =32'b00000000000000000000000000000000;
8'b10000011 : Out =32'b00000000000000000000000000000000;
8'b10000100 : Out =32'b00000000000000000000000000000000;
8'b10000101 : Out =32'b00000000000000000000000000000000;
8'b10000110 : Out =32'b00000000000000000000000000000000;
8'b10000111 : Out =32'b00000000000000000000000000000000;
8'b10001000 : Out =32'b00000000000000000000000000000000;
8'b10001001 : Out =32'b00000000000000000000000000000000;
8'b10001010 : Out =32'b00000000000000000000000000000000;
8'b10001011 : Out =32'b00000000000000000000000000000000;
8'b10001100 : Out =32'b00000000000000000000000000000000;
8'b10001101 : Out =32'b00000000000000000000000000000000;
8'b10001110 : Out =32'b00000000000000000000000000000000;
8'b10001111 : Out =32'b00000000000000000000000000000000;
8'b10010000 : Out =32'b00000000000000000000000000000000;
8'b10010001 : Out =32'b00000000000000000000000000000000;
8'b10010010 : Out =32'b00000000000000000000000000000000;
8'b10010011 : Out =32'b00000000000000000000000000000000;
8'b10010100 : Out =32'b00000000000000000000000000000000;
8'b10010101 : Out =32'b00000000000000000000000000000000;
8'b10010110 : Out =32'b00000000000000000000000000000000;
8'b10010111 : Out =32'b00000000000000000000000000000000;
8'b10011000 : Out =32'b00000000000000000000000000000000;
8'b10011001 : Out =32'b00000000000000000000000000000000;
8'b10011010 : Out =32'b00000000000000000000000000000000;
8'b10011011 : Out =32'b00000000000000000000000000000000;
8'b10011100 : Out =32'b00000000000000000000000000000000;
8'b10011101 : Out =32'b00000000000000000000000000000000;
8'b10011110 : Out =32'b00000000000000000000000000000000;
8'b10011111 : Out =32'b00000000000000000000000000000000;
8'b10100000 : Out =32'b00000000000000000000000000000000;
8'b10100001 : Out =32'b00000000000000000000000000000000;
8'b10100010 : Out =32'b00000000000000000000000000000000;
8'b10100011 : Out =32'b00000000000000000000000000000000;
8'b10100100 : Out =32'b00000000000000000000000000000000;
8'b10100101 : Out =32'b00000000000000000000000000000001;
8'b10100110 : Out =32'b00000000000000000000000000000001;
8'b10100111 : Out =32'b00000000000000000000000000000001;
8'b10101000 : Out =32'b00000000000000000000000000000001;
8'b10101001 : Out =32'b00000000000000000000000000000010;
8'b10101010 : Out =32'b00000000000000000000000000000010;
8'b10101011 : Out =32'b00000000000000000000000000000011;
8'b10101100 : Out =32'b00000000000000000000000000000011;
8'b10101101 : Out =32'b00000000000000000000000000000100;
8'b10101110 : Out =32'b00000000000000000000000000000101;
8'b10101111 : Out =32'b00000000000000000000000000000111;
8'b10110000 : Out =32'b00000000000000000000000000001001;
8'b10110001 : Out =32'b00000000000000000000000000001011;
8'b10110010 : Out =32'b00000000000000000000000000001111;
8'b10110011 : Out =32'b00000000000000000000000000010011;
8'b10110100 : Out =32'b00000000000000000000000000011000;
8'b10110101 : Out =32'b00000000000000000000000000011111;
8'b10110110 : Out =32'b00000000000000000000000000101000;
8'b10110111 : Out =32'b00000000000000000000000000110011;
8'b10111000 : Out =32'b00000000000000000000000001000001;
8'b10111001 : Out =32'b00000000000000000000000001010100;
8'b10111010 : Out =32'b00000000000000000000000001101100;
8'b10111011 : Out =32'b00000000000000000000000010001010;
8'b10111100 : Out =32'b00000000000000000000000010110010;
8'b10111101 : Out =32'b00000000000000000000000011100100;
8'b10111110 : Out =32'b00000000000000000000000100100101;
8'b10111111 : Out =32'b00000000000000000000000101111000;
8'b11000000 : Out =32'b00000000000000000000000111100011;
8'b11000001 : Out =32'b00000000000000000000001001101101;
8'b11000010 : Out =32'b00000000000000000000001100011101;
8'b11000011 : Out =32'b00000000000000000000001111111111;
8'b11000100 : Out =32'b00000000000000000000010100100010;
8'b11000101 : Out =32'b00000000000000000000011010010111;
8'b11000110 : Out =32'b00000000000000000000100001110110;
8'b11000111 : Out =32'b00000000000000000000101011011101;
8'b11001000 : Out =32'b00000000000000000000110111110011;
8'b11001001 : Out =32'b00000000000000000001000111101010;
8'b11001010 : Out =32'b00000000000000000001011100000000;
8'b11001011 : Out =32'b00000000000000000001110110001001;
8'b11001100 : Out =32'b00000000000000000010010111101100;
8'b11001101 : Out =32'b00000000000000000011000010110001;
8'b11001110 : Out =32'b00000000000000000011111010000110;
8'b11001111 : Out =32'b00000000000000000101000001001000;
8'b11010000 : Out =32'b00000000000000000110011100010101;
8'b11010001 : Out =32'b00000000000000001000010001011100;
8'b11010010 : Out =32'b00000000000000001010100111110100;
8'b11010011 : Out =32'b00000000000000001101101000111001;
8'b11010100 : Out =32'b00000000000000010001100000110100;
8'b11010101 : Out =32'b00000000000000010110011111001001;
8'b11010110 : Out =32'b00000000000000011100110111111001;
8'b11010111 : Out =32'b00000000000000100101000100101110;
8'b11011000 : Out =32'b00000000000000101111100110100110;
8'b11011001 : Out =32'b00000000000000111101000111110111;
8'b11011010 : Out =32'b00000000000001001110011110110110;
8'b11011011 : Out =32'b00000000000001100100110001010101;
8'b11011100 : Out =32'b00000000000010000001011000111000;
8'b11011101 : Out =32'b00000000000010100110001000011110;
8'b11011110 : Out =32'b00000000000011010101010011110000;
8'b11011111 : Out =32'b00000000000100010001111000001100;
8'b11100000 : Out =32'b00000000000101011111101000111110;
8'b11100001 : Out =32'b00000000000111000011011110001101;
8'b11100010 : Out =32'b00000000001001000011101000010110;
8'b11100011 : Out =32'b00000000001011101000001001001011;
8'b11100100 : Out =32'b00000000001110111011010011100111;
8'b11100101 : Out =32'b00000000010011001010010100100000;
8'b11100110 : Out =32'b00000000011000100110000110101001;
8'b11100111 : Out =32'b00000000011111100100010100111110;
8'b11101000 : Out =32'b00000000101000100000101110111100;
8'b11101001 : Out =32'b00000000110011111110110011001001;
8'b11101010 : Out =32'b00000001000010101011110110010100;
8'b11101011 : Out =32'b00000001010101100001101100101101;
8'b11101100 : Out =32'b00000001101101101001111101101000;
8'b11101101 : Out =32'b00000010001100100010001001010011;
8'b11101110 : Out =32'b00000010110100000000101001001111;
8'b11101111 : Out =32'b00000011100110011010110010000010;
8'b11110000 : Out =32'b00000100100110101011111010001000;
8'b11110001 : Out =32'b00000101111000011101100001001100;
8'b11110010 : Out =32'b00000111100000010000000110100000;
8'b11110011 : Out =32'b00001001100011100100000101000000;
8'b11110100 : Out =32'b00001100001001000001101000011110;
8'b11110101 : Out =32'b00001111011000011101011010110101;
8'b11110110 : Out =32'b00010011011010110111000100010010;
8'b11110111 : Out =32'b00011000011010001101001010010001;
8'b11111000 : Out =32'b00011110100001000001010100101100;
8'b11111001 : Out =32'b00100101111001100110101111010010;
8'b11111010 : Out =32'b00101110101100110111000001101011;
8'b11111011 : Out =32'b00111001000000101110000001010101;
8'b11111100 : Out =32'b01000100110110010101100001010001;
8'b11111101 : Out =32'b01010010001000010101100001000011;
8'b11111110 : Out =32'b01100000101001101000000101011001;
8'b11111111 : Out =32'b01110000000101010011001101101010;
8'b00000000 : Out =32'b10000000000000000000000000000000;
8'b00000001 : Out =32'b10001111111010101100110010010110;
8'b00000010 : Out =32'b10011111010110010111111010100111;
8'b00000011 : Out =32'b10101101110111101010011110111101;
8'b00000100 : Out =32'b10111011001001101010011110101111;
8'b00000101 : Out =32'b11000110111111010001111110101011;
8'b00000110 : Out =32'b11010001010011001000111110010101;
8'b00000111 : Out =32'b11011010000110011001010000101110;
8'b00001000 : Out =32'b11100001011110111110101011010100;
8'b00001001 : Out =32'b11100111100101110010110101101111;
8'b00001010 : Out =32'b11101100100101001000111011101110;
8'b00001011 : Out =32'b11110000100111100010100101001011;
8'b00001100 : Out =32'b11110011110110111110010111100010;
8'b00001101 : Out =32'b11110110011100011011111011000000;
8'b00001110 : Out =32'b11111000011111101111111001100000;
8'b00001111 : Out =32'b11111010000111100010011110110100;
8'b00010000 : Out =32'b11111011011001010100000101111000;
8'b00010001 : Out =32'b11111100011001100101001101111110;
8'b00010010 : Out =32'b11111101001011111111010110110001;
8'b00010011 : Out =32'b11111101110011011101110110101101;
8'b00010100 : Out =32'b11111110010010010110000010011000;
8'b00010101 : Out =32'b11111110101010011110010011010011;
8'b00010110 : Out =32'b11111110111101010100001001101100;
8'b00010111 : Out =32'b11111111001100000001001100110111;
8'b00011000 : Out =32'b11111111010111011111010001000100;
8'b00011001 : Out =32'b11111111100000011011101011000010;
8'b00011010 : Out =32'b11111111100111011001111001010111;
8'b00011011 : Out =32'b11111111101100110101101011100000;
8'b00011100 : Out =32'b11111111110001000100101100011001;
8'b00011101 : Out =32'b11111111110100010111110110110101;
8'b00011110 : Out =32'b11111111110110111100010111101010;
8'b00011111 : Out =32'b11111111111000111100100001110011;
8'b00100000 : Out =32'b11111111111010100000010111000010;
8'b00100001 : Out =32'b11111111111011101110000111110100;
8'b00100010 : Out =32'b11111111111100101010101100010000;
8'b00100011 : Out =32'b11111111111101011001110111100010;
8'b00100100 : Out =32'b11111111111101111110100111001000;
8'b00100101 : Out =32'b11111111111110011011001110101011;
8'b00100110 : Out =32'b11111111111110110001100001001010;
8'b00100111 : Out =32'b11111111111111000010111000001001;
8'b00101000 : Out =32'b11111111111111010000011001011010;
8'b00101001 : Out =32'b11111111111111011010111011010010;
8'b00101010 : Out =32'b11111111111111100011001000000111;
8'b00101011 : Out =32'b11111111111111101001100000110111;
8'b00101100 : Out =32'b11111111111111101110011111001100;
8'b00101101 : Out =32'b11111111111111110010010111000111;
8'b00101110 : Out =32'b11111111111111110101011000001100;
8'b00101111 : Out =32'b11111111111111110111101110100100;
8'b00110000 : Out =32'b11111111111111111001100011101011;
8'b00110001 : Out =32'b11111111111111111010111110111000;
8'b00110010 : Out =32'b11111111111111111100000101111010;
8'b00110011 : Out =32'b11111111111111111100111101001111;
8'b00110100 : Out =32'b11111111111111111101101000010100;
8'b00110101 : Out =32'b11111111111111111110001001110111;
8'b00110110 : Out =32'b11111111111111111110100100000000;
8'b00110111 : Out =32'b11111111111111111110111000010110;
8'b00111000 : Out =32'b11111111111111111111001000001101;
8'b00111001 : Out =32'b11111111111111111111010100100011;
8'b00111010 : Out =32'b11111111111111111111011110001010;
8'b00111011 : Out =32'b11111111111111111111100101101001;
8'b00111100 : Out =32'b11111111111111111111101011011110;
8'b00111101 : Out =32'b11111111111111111111110000000001;
8'b00111110 : Out =32'b11111111111111111111110011100011;
8'b00111111 : Out =32'b11111111111111111111110110010011;
8'b01000000 : Out =32'b11111111111111111111111000011101;
8'b01000001 : Out =32'b11111111111111111111111010001000;
8'b01000010 : Out =32'b11111111111111111111111011011011;
8'b01000011 : Out =32'b11111111111111111111111100011100;
8'b01000100 : Out =32'b11111111111111111111111101001110;
8'b01000101 : Out =32'b11111111111111111111111101110110;
8'b01000110 : Out =32'b11111111111111111111111110010100;
8'b01000111 : Out =32'b11111111111111111111111110101100;
8'b01001000 : Out =32'b11111111111111111111111110111111;
8'b01001001 : Out =32'b11111111111111111111111111001101;
8'b01001010 : Out =32'b11111111111111111111111111011000;
8'b01001011 : Out =32'b11111111111111111111111111100001;
8'b01001100 : Out =32'b11111111111111111111111111101000;
8'b01001101 : Out =32'b11111111111111111111111111101101;
8'b01001110 : Out =32'b11111111111111111111111111110001;
8'b01001111 : Out =32'b11111111111111111111111111110101;
8'b01010000 : Out =32'b11111111111111111111111111110111;
8'b01010001 : Out =32'b11111111111111111111111111111001;
8'b01010010 : Out =32'b11111111111111111111111111111011;
8'b01010011 : Out =32'b11111111111111111111111111111100;
8'b01010100 : Out =32'b11111111111111111111111111111101;
8'b01010101 : Out =32'b11111111111111111111111111111101;
8'b01010110 : Out =32'b11111111111111111111111111111110;
8'b01010111 : Out =32'b11111111111111111111111111111110;
8'b01011000 : Out =32'b11111111111111111111111111111111;
8'b01011001 : Out =32'b11111111111111111111111111111111;
8'b01011010 : Out =32'b11111111111111111111111111111111;
8'b01011011 : Out =32'b11111111111111111111111111111111;
8'b01011100 : Out =32'b11111111111111111111111111111111;
8'b01011101 : Out =32'b11111111111111111111111111111111;
8'b01011110 : Out =32'b11111111111111111111111111111111;
8'b01011111 : Out =32'b11111111111111111111111111111111;
8'b01100000 : Out =32'b11111111111111111111111111111111;
8'b01100001 : Out =32'b11111111111111111111111111111111;
8'b01100010 : Out =32'b11111111111111111111111111111111;
8'b01100011 : Out =32'b11111111111111111111111111111111;
8'b01100100 : Out =32'b11111111111111111111111111111111;
8'b01100101 : Out =32'b11111111111111111111111111111111;
8'b01100110 : Out =32'b11111111111111111111111111111111;
8'b01100111 : Out =32'b11111111111111111111111111111111;
8'b01101000 : Out =32'b11111111111111111111111111111111;
8'b01101001 : Out =32'b11111111111111111111111111111111;
8'b01101010 : Out =32'b11111111111111111111111111111111;
8'b01101011 : Out =32'b11111111111111111111111111111111;
8'b01101100 : Out =32'b11111111111111111111111111111111;
8'b01101101 : Out =32'b11111111111111111111111111111111;
8'b01101110 : Out =32'b11111111111111111111111111111111;
8'b01101111 : Out =32'b11111111111111111111111111111111;
8'b01110000 : Out =32'b11111111111111111111111111111111;
8'b01110001 : Out =32'b11111111111111111111111111111111;
8'b01110010 : Out =32'b11111111111111111111111111111111;
8'b01110011 : Out =32'b11111111111111111111111111111111;
8'b01110100 : Out =32'b11111111111111111111111111111111;
8'b01110101 : Out =32'b11111111111111111111111111111111;
8'b01110110 : Out =32'b11111111111111111111111111111111;
8'b01110111 : Out =32'b11111111111111111111111111111111;
8'b01111000 : Out =32'b11111111111111111111111111111111;
8'b01111001 : Out =32'b11111111111111111111111111111111;
8'b01111010 : Out =32'b11111111111111111111111111111111;
8'b01111011 : Out =32'b11111111111111111111111111111111;
8'b01111100 : Out =32'b11111111111111111111111111111111;
8'b01111101 : Out =32'b11111111111111111111111111111111;
8'b01111110 : Out =32'b11111111111111111111111111111111;
8'b01111111 : Out =32'b11111111111111111111111111111111;

endcase
end
endmodule